`timescale 1ns / 10ps

module tb();
	reg CLK;
	initial begin
		CLK = 1'b0;
		forever #5 CLK = ~CLK;
	end
	
	reg [15:0] OP1_i, OP2_i;
	wire [15:0] MUL_o;
	FPMUL umul (OP1_i, OP2_i, MUL_o);
	initial begin
		OP1_i = 16'b0100000110000000; OP2_i = 16'b0011101000000000; // 2.75, 0.75
        #(10) OP1_i = 16'b0100000000000000; OP2_i = 16'b0011111000000000; 
        #(10) OP1_i = 16'b0111100011000000; OP2_i = 16'b0111011100000100;	//overflow
        #(10) OP1_i = 16'b0000100000000000; OP2_i = 16'b0001011100000000;	//underflow
		#(10) OP1_i = 16'b0000000000000000; OP2_i = 16'b0000000000000000;	//underflow
		#(10) OP1_i = 16'b0100001001001001; OP2_i = 16'b1100001001100110;	
		#(10) OP1_i = 16'b0011110100000000; OP2_i = 16'b0011110100000000; 
		#(10) OP1_i = 16'b0011111000000000; OP2_i = 16'b0011111000000000; 
		#(10) OP1_i = 16'b0011111110000000; OP2_i = 16'b0011111110000000; 
		#(10) OP1_i = 16'b0101110100000000; OP2_i = 16'b0101110100000000; //overflow
		#(10) OP1_i = 16'b0101101000000000; OP2_i = 16'b0101111000000000; //overflow 
		#(10) OP1_i = 16'b0101101110000000; OP2_i = 16'b0101111110000000; //overflow 
		#(10) OP1_i = 16'b0010000100000000; OP2_i = 16'b0001110100000000; //underflow 
		#(10) OP1_i = 16'b0001111000000000; OP2_i = 16'b0001111000000000; //underflow
		#(10) OP1_i = 16'b0001111000000000; OP2_i = 16'b0010001000000000; 
		#(10) OP1_i = 16'b0001111110000000; OP2_i = 16'b0001111110000000; //underflow
		#(10) OP1_i = 16'b0001111110000000; OP2_i = 16'b0010001110000000; 
		#(20)
		$finish();
	end	

	initial begin
		$dumpfile("fpmultest.dmp");
		$dumpvars;
	end

endmodule
	/*
		//차재민 tb	
		OP1_i = 16'b0011110100000000; OP2_i = 16'b0011110100000000; //normalized 0011111001000000
		#(10) OP1_i = 16'b0011111000000000; OP2_i = 16'b0011111000000000; //normal 0100000010000000
		#(10) OP1_i = 16'b0011111110000000; OP2_i = 16'b0011111110000000; //normal 0100001100001000
		#(10) OP1_i = 16'b0101110100000000; OP2_i = 16'b0101110100000000; //(1.01 2^8 * 1.01 2^8) 오버플로우 0111110000000000
		#(10) OP1_i = 16'b0101101000000000; OP2_i = 16'b0101111000000000; //(1.1 2^7 * 1.1 2^8) 오버플로우 0111110000000000
		#(10) OP1_i = 16'b0101101110000000; OP2_i = 16'b0101111110000000; //(1.111 2^7 * 1.111 2^8) 오버플로우 0111110000000000
		#(10) OP1_i = 16'b0010000100000000; OP2_i = 16'b0001110100000000; //(1.01 2^-7 * 1.01 2^-8) 언더플로우 0000000000000000
		#(10) OP1_i = 16'b0001111000000000; OP2_i = 16'b0001111000000000; //(1.1 2^-8 * 1.1 2^-8) 언더플로우 0000000000000000
		#(10) OP1_i = 16'b0001111000000000; OP2_i = 16'b0010001000000000; //(1.1 2^-8 * 1.1 2^-7) normal 0000010010000000
		#(10) OP1_i = 16'b0001111110000000; OP2_i = 16'b0001111110000000; //(1.111 2^-8 * 1.111 2^-8) 언더플로우 0000000000000000
		#(10) OP1_i = 16'b0001111110000000; OP2_i = 16'b0010001110000000; //(1.111 2^-8 * 1.111 2^-7) normal 0000011100001000
	*/