`timescale 1ns / 10ps

module tb();

	reg CLK;

	initial begin
		CLK = 1'b0;
		forever #5 CLK = ~CLK;
	end
	
	reg [15:0] OP1_i, OP2_i;
	wire [15:0] ADD_o;

	FPADD uadd (OP1_i, OP2_i, ADD_o);

	initial begin
		/*
		OP1_i = 16'b0011110001100000; OP2_i = 16'b0011110000000000; 
        #(10) OP1_i = 16'b0010000001100000; OP2_i = 16'b0011110100000000;
		#(10) OP1_i = 16'b0011110001100000; OP2_i = 16'b0011110000000000; 
		#(10) OP1_i = 16'b0011110001100000; OP2_i = 16'b1011110000000000; 
		#(10) OP1_i = 16'b0011110001100000; OP2_i = 16'b0011110000000000; 0100000000110000
		#(10) OP1_i = 16'b0011110001100000; OP2_i = 16'b1011110000000000; //0010111000000000
		#(10) OP1_i = 16'b0010000001100000; OP2_i = 16'b0011110100000000; //0011110100001000
		#(10) OP1_i = 16'b0100000000000000; OP2_i = 16'b0100010000000000; //0100011000000000
		#(10) OP1_i = 16'b0100010000100000; OP2_i = 16'b1100010000000000; //0011000000000000
		
		//underflow
		#(10) OP1_i = 16'b0000010000100000; OP2_i = 16'b1000000000000010; //0000000000000000
		
		//overflow
		#(10) OP1_i = 16'b0111101000000000; OP2_i = 16'b0111011000000000; //0111110000000000
		#(10) OP1_i = 16'b0111101000000000; OP2_i = 16'b0111101000000000;
		*/
		
		//(+)+(+)
		OP1_i = 16'b0101000000000000; OP2_i = 16'b0101000000000000; //0101010000000000
		#(10) OP1_i = 16'b0101001100000000; OP2_i = 16'b0101001100000000; //0101011100000000 
		#(10) OP1_i = 16'b0100100000000000; OP2_i = 16'b0101100000000000; //0101100001000000 
		#(10) OP1_i = 16'b0100101100000000; OP2_i = 16'b0101101111000000; //0101110000011000 
		#(10) OP1_i = 16'b0000100000000000; OP2_i = 16'b0000100000000000; //0000110000000000 
		#(10) OP1_i = 16'b0000111100000000; OP2_i = 16'b0101101100000000; //0101101100000000 
		#(10) OP1_i = 16'b0011001100000000; OP2_i = 16'b0100001100000000; //0100001101110000 
		//overflow
		#(10) OP1_i = 16'b0111100000000000; OP2_i = 16'b0111100000000000; //0111110000000000 
		#(10) OP1_i = 16'b0111011100000000; OP2_i = 16'b0111101110000000; //0111110000000000 
		#(10) OP1_i = 16'b0111101111111111; OP2_i = 16'b0101000000000000; //0111110000000000 
		//(-)+(-)
		#(10) OP1_i = 16'b1101001100000000; OP2_i = 16'b1101001100000000; //1101011100000000 
		#(10) OP1_i = 16'b1100100000000000; OP2_i = 16'b1101100000000000; //1101100001000000 
		#(10) OP1_i = 16'b1100101100000000; OP2_i = 16'b1101101111000000; //1101110000011000 
		#(10) OP1_i = 16'b1000100000000000; OP2_i = 16'b1000100000000000; //1000110000000000 
		#(10) OP1_i = 16'b1000111100000000; OP2_i = 16'b1101101100000000; //1101101100000000 
		#(10) OP1_i = 16'b1011001100000000; OP2_i = 16'b1100001100000000; //1100001101110000 
		//(-)overflow
		#(10) OP1_i = 16'b1111100000000000; OP2_i = 16'b1111100000000000; //1111110000000000 
		#(10) OP1_i = 16'b1111011100000000; OP2_i = 16'b1111101110000000; //1111110000000000 
		#(10) OP1_i = 16'b1111101111111111; OP2_i = 16'b1101000000000000; //1111110000000000 
		//(+)+(-)
		#(10) OP1_i = 16'b0100110000000001; OP2_i = 16'b1100100000000000; //0100100000000010 
		#(10) OP1_i = 16'b0100111111111111; OP2_i = 16'b1100100000000000; //0100110111111111 
		#(10) OP1_i = 16'b0101000000000000; OP2_i = 16'b1100000000000000; //0100111110000000 
		#(10) OP1_i = 16'b0101001111111111; OP2_i = 16'b1100001111111111; //0101001110000000 
		#(10) OP1_i = 16'b0101010000000000; OP2_i = 16'b1100111111111111; //0101000000000010 
		#(10) OP1_i = 16'b0101011111111110; OP2_i = 16'b1100111111111111; //0101010111111111 
		#(10) OP1_i = 16'b0101001111111111; OP2_i = 16'b1101000000000000; //0100111111111110 
		//same exp
		#(10) OP1_i = 16'b0100011111111111; OP2_i = 16'b1100011111111111; //0000000000000000 
		#(10) OP1_i = 16'b0101010000000000; OP2_i = 16'b1101011111111111; //1101001111111110 
		//(+)+(-)
		#(10) OP1_i = 16'b0100111111111111; OP2_i = 16'b1101001111111110; //1100111111111110 
		#(10) OP1_i = 16'b0100101111111111; OP2_i = 16'b1101001111111110; //1101000111111111 
		#(10) OP1_i = 16'b0100110000000000; OP2_i = 16'b1101010000000000; //1101001000000000 
		#(10) OP1_i = 16'b0100011111111111; OP2_i = 16'b1101011111111111; //1101011110000000 
		#(10) OP1_i = 16'b0100000000000000; OP2_i = 16'b1101000000000001; //1100111110000010 
		#(10) OP1_i = 16'b0100000000000000; OP2_i = 16'b1100111111111111; //1100111101111111 
		//underflow
		#(10) OP1_i = 16'b0000100000000000; OP2_i = 16'b1000011111111111; //0000000000000000
		#(10) OP1_i = 16'b0000011111111111; OP2_i = 16'b1000011111111110; //0000000000000000
		#(10) OP1_i = 16'b0000010000000000; OP2_i = 16'b1000010000000001; //0000000000000000 
		//input oveflow/0
		#(10) OP1_i = 16'b0111110000000000; OP2_i = 16'b1010110000100001; //1111110000000000
		#(10) OP1_i = 16'b0000000000000000; OP2_i = 16'b0001000000100001; //0111110000000000
        #(10) OP1_i=0; OP2_i=0;	//0000000000000000
		#(20)
		
		$finish();
	end


	initial begin
		$dumpfile("fpaddtest.dmp");
		$dumpvars;
	end

endmodule



